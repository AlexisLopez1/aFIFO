package tb_fifo_pkg;
    localparam DW = 8;
    typedef logic [DW-1:0]  data_t;
endpackage